VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mprj_logic_high
  CLASS BLOCK ;
  FOREIGN mprj_logic_high ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 23.000 ;
  PIN HI[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 19.000 165.050 23.000 ;
    END
  END HI[0]
  PIN HI[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 9.560 300.000 10.160 ;
    END
  END HI[100]
  PIN HI[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 19.000 144.810 23.000 ;
    END
  END HI[101]
  PIN HI[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END HI[102]
  PIN HI[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END HI[103]
  PIN HI[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 19.000 47.290 23.000 ;
    END
  END HI[104]
  PIN HI[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END HI[105]
  PIN HI[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END HI[106]
  PIN HI[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 19.000 102.490 23.000 ;
    END
  END HI[107]
  PIN HI[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END HI[108]
  PIN HI[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 19.000 65.690 23.000 ;
    END
  END HI[109]
  PIN HI[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END HI[10]
  PIN HI[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END HI[110]
  PIN HI[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 19.000 258.890 23.000 ;
    END
  END HI[111]
  PIN HI[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END HI[112]
  PIN HI[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 19.000 141.130 23.000 ;
    END
  END HI[113]
  PIN HI[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END HI[114]
  PIN HI[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END HI[115]
  PIN HI[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END HI[116]
  PIN HI[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 19.000 95.130 23.000 ;
    END
  END HI[117]
  PIN HI[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 19.000 234.970 23.000 ;
    END
  END HI[118]
  PIN HI[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END HI[119]
  PIN HI[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 19.000 191.730 23.000 ;
    END
  END HI[11]
  PIN HI[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END HI[120]
  PIN HI[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 19.000 63.850 23.000 ;
    END
  END HI[121]
  PIN HI[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 19.000 51.890 23.000 ;
    END
  END HI[122]
  PIN HI[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 19.000 74.890 23.000 ;
    END
  END HI[123]
  PIN HI[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 19.000 59.250 23.000 ;
    END
  END HI[124]
  PIN HI[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END HI[125]
  PIN HI[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 19.000 231.290 23.000 ;
    END
  END HI[126]
  PIN HI[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 19.000 188.970 23.000 ;
    END
  END HI[127]
  PIN HI[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 19.000 272.690 23.000 ;
    END
  END HI[128]
  PIN HI[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END HI[129]
  PIN HI[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END HI[12]
  PIN HI[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 19.000 200.930 23.000 ;
    END
  END HI[130]
  PIN HI[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 19.000 98.810 23.000 ;
    END
  END HI[131]
  PIN HI[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END HI[132]
  PIN HI[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 19.000 18.770 23.000 ;
    END
  END HI[133]
  PIN HI[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 19.000 273.610 23.000 ;
    END
  END HI[134]
  PIN HI[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 19.000 216.570 23.000 ;
    END
  END HI[135]
  PIN HI[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 19.000 292.010 23.000 ;
    END
  END HI[136]
  PIN HI[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 19.000 66.610 23.000 ;
    END
  END HI[137]
  PIN HI[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 19.000 21.530 23.000 ;
    END
  END HI[138]
  PIN HI[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END HI[139]
  PIN HI[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END HI[13]
  PIN HI[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 19.000 194.490 23.000 ;
    END
  END HI[140]
  PIN HI[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 19.000 294.770 23.000 ;
    END
  END HI[141]
  PIN HI[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END HI[142]
  PIN HI[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END HI[143]
  PIN HI[144]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 19.000 30.730 23.000 ;
    END
  END HI[144]
  PIN HI[145]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 19.000 219.330 23.000 ;
    END
  END HI[145]
  PIN HI[146]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 19.000 131.930 23.000 ;
    END
  END HI[146]
  PIN HI[147]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 19.000 296.610 23.000 ;
    END
  END HI[147]
  PIN HI[148]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 19.000 96.050 23.000 ;
    END
  END HI[148]
  PIN HI[149]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END HI[149]
  PIN HI[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END HI[14]
  PIN HI[150]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END HI[150]
  PIN HI[151]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 19.000 198.170 23.000 ;
    END
  END HI[151]
  PIN HI[152]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 19.000 174.250 23.000 ;
    END
  END HI[152]
  PIN HI[153]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END HI[153]
  PIN HI[154]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 19.000 93.290 23.000 ;
    END
  END HI[154]
  PIN HI[155]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 19.000 261.650 23.000 ;
    END
  END HI[155]
  PIN HI[156]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END HI[156]
  PIN HI[157]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END HI[157]
  PIN HI[158]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END HI[158]
  PIN HI[159]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END HI[159]
  PIN HI[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END HI[15]
  PIN HI[160]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END HI[160]
  PIN HI[161]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 19.000 267.170 23.000 ;
    END
  END HI[161]
  PIN HI[162]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 19.000 221.170 23.000 ;
    END
  END HI[162]
  PIN HI[163]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 19.000 185.290 23.000 ;
    END
  END HI[163]
  PIN HI[164]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 19.000 39.010 23.000 ;
    END
  END HI[164]
  PIN HI[165]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 19.000 195.410 23.000 ;
    END
  END HI[165]
  PIN HI[166]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END HI[166]
  PIN HI[167]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 19.000 153.090 23.000 ;
    END
  END HI[167]
  PIN HI[168]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END HI[168]
  PIN HI[169]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 19.000 26.130 23.000 ;
    END
  END HI[169]
  PIN HI[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 19.000 15.090 23.000 ;
    END
  END HI[16]
  PIN HI[170]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END HI[170]
  PIN HI[171]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END HI[171]
  PIN HI[172]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END HI[172]
  PIN HI[173]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 19.000 278.210 23.000 ;
    END
  END HI[173]
  PIN HI[174]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 19.000 212.890 23.000 ;
    END
  END HI[174]
  PIN HI[175]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END HI[175]
  PIN HI[176]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END HI[176]
  PIN HI[177]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END HI[177]
  PIN HI[178]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 19.000 108.010 23.000 ;
    END
  END HI[178]
  PIN HI[179]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 19.000 165.970 23.000 ;
    END
  END HI[179]
  PIN HI[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END HI[17]
  PIN HI[180]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END HI[180]
  PIN HI[181]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END HI[181]
  PIN HI[182]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END HI[182]
  PIN HI[183]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 19.000 263.490 23.000 ;
    END
  END HI[183]
  PIN HI[184]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 19.000 123.650 23.000 ;
    END
  END HI[184]
  PIN HI[185]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END HI[185]
  PIN HI[186]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 19.000 27.050 23.000 ;
    END
  END HI[186]
  PIN HI[187]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END HI[187]
  PIN HI[188]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 19.000 177.930 23.000 ;
    END
  END HI[188]
  PIN HI[189]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 19.000 206.450 23.000 ;
    END
  END HI[189]
  PIN HI[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 19.000 72.130 23.000 ;
    END
  END HI[18]
  PIN HI[190]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END HI[190]
  PIN HI[191]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 19.000 113.530 23.000 ;
    END
  END HI[191]
  PIN HI[192]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 19.000 62.930 23.000 ;
    END
  END HI[192]
  PIN HI[193]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 19.000 8.650 23.000 ;
    END
  END HI[193]
  PIN HI[194]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END HI[194]
  PIN HI[195]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END HI[195]
  PIN HI[196]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 19.000 209.210 23.000 ;
    END
  END HI[196]
  PIN HI[197]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 19.000 117.210 23.000 ;
    END
  END HI[197]
  PIN HI[198]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END HI[198]
  PIN HI[199]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END HI[199]
  PIN HI[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 19.000 158.610 23.000 ;
    END
  END HI[19]
  PIN HI[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END HI[1]
  PIN HI[200]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END HI[200]
  PIN HI[201]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END HI[201]
  PIN HI[202]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END HI[202]
  PIN HI[203]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END HI[203]
  PIN HI[204]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END HI[204]
  PIN HI[205]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 19.000 39.930 23.000 ;
    END
  END HI[205]
  PIN HI[206]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 19.000 170.570 23.000 ;
    END
  END HI[206]
  PIN HI[207]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 19.000 120.890 23.000 ;
    END
  END HI[207]
  PIN HI[208]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END HI[208]
  PIN HI[209]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END HI[209]
  PIN HI[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END HI[20]
  PIN HI[210]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 19.000 183.450 23.000 ;
    END
  END HI[210]
  PIN HI[211]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END HI[211]
  PIN HI[212]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END HI[212]
  PIN HI[213]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END HI[213]
  PIN HI[214]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END HI[214]
  PIN HI[215]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END HI[215]
  PIN HI[216]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END HI[216]
  PIN HI[217]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 19.000 42.690 23.000 ;
    END
  END HI[217]
  PIN HI[218]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 19.000 276.370 23.000 ;
    END
  END HI[218]
  PIN HI[219]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END HI[219]
  PIN HI[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 19.000 138.370 23.000 ;
    END
  END HI[21]
  PIN HI[220]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END HI[220]
  PIN HI[221]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END HI[221]
  PIN HI[222]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END HI[222]
  PIN HI[223]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END HI[223]
  PIN HI[224]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 19.000 222.090 23.000 ;
    END
  END HI[224]
  PIN HI[225]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 19.000 4.050 23.000 ;
    END
  END HI[225]
  PIN HI[226]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 15.000 300.000 15.600 ;
    END
  END HI[226]
  PIN HI[227]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 19.000 254.290 23.000 ;
    END
  END HI[227]
  PIN HI[228]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END HI[228]
  PIN HI[229]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 19.000 236.810 23.000 ;
    END
  END HI[229]
  PIN HI[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END HI[22]
  PIN HI[230]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 19.000 197.250 23.000 ;
    END
  END HI[230]
  PIN HI[231]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END HI[231]
  PIN HI[232]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END HI[232]
  PIN HI[233]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 19.000 57.410 23.000 ;
    END
  END HI[233]
  PIN HI[234]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END HI[234]
  PIN HI[235]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END HI[235]
  PIN HI[236]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 19.000 23.370 23.000 ;
    END
  END HI[236]
  PIN HI[237]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END HI[237]
  PIN HI[238]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 19.000 156.770 23.000 ;
    END
  END HI[238]
  PIN HI[239]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END HI[239]
  PIN HI[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END HI[23]
  PIN HI[240]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END HI[240]
  PIN HI[241]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 19.000 211.050 23.000 ;
    END
  END HI[241]
  PIN HI[242]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 19.000 281.890 23.000 ;
    END
  END HI[242]
  PIN HI[243]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 19.000 255.210 23.000 ;
    END
  END HI[243]
  PIN HI[244]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 19.000 45.450 23.000 ;
    END
  END HI[244]
  PIN HI[245]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END HI[245]
  PIN HI[246]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END HI[246]
  PIN HI[247]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 19.000 36.250 23.000 ;
    END
  END HI[247]
  PIN HI[248]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 19.000 85.010 23.000 ;
    END
  END HI[248]
  PIN HI[249]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END HI[249]
  PIN HI[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 19.000 207.370 23.000 ;
    END
  END HI[24]
  PIN HI[250]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 17.720 300.000 18.320 ;
    END
  END HI[250]
  PIN HI[251]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END HI[251]
  PIN HI[252]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 19.000 239.570 23.000 ;
    END
  END HI[252]
  PIN HI[253]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 19.000 128.250 23.000 ;
    END
  END HI[253]
  PIN HI[254]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END HI[254]
  PIN HI[255]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END HI[255]
  PIN HI[256]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 19.000 227.610 23.000 ;
    END
  END HI[256]
  PIN HI[257]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 19.000 246.930 23.000 ;
    END
  END HI[257]
  PIN HI[258]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END HI[258]
  PIN HI[259]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 19.000 61.090 23.000 ;
    END
  END HI[259]
  PIN HI[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 19.000 108.930 23.000 ;
    END
  END HI[25]
  PIN HI[260]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 19.000 149.410 23.000 ;
    END
  END HI[260]
  PIN HI[261]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END HI[261]
  PIN HI[262]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END HI[262]
  PIN HI[263]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 19.000 111.690 23.000 ;
    END
  END HI[263]
  PIN HI[264]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END HI[264]
  PIN HI[265]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END HI[265]
  PIN HI[266]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END HI[266]
  PIN HI[267]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 19.000 130.090 23.000 ;
    END
  END HI[267]
  PIN HI[268]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END HI[268]
  PIN HI[269]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 19.000 243.250 23.000 ;
    END
  END HI[269]
  PIN HI[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END HI[26]
  PIN HI[270]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END HI[270]
  PIN HI[271]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 19.000 284.650 23.000 ;
    END
  END HI[271]
  PIN HI[272]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 19.000 137.450 23.000 ;
    END
  END HI[272]
  PIN HI[273]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 19.000 186.210 23.000 ;
    END
  END HI[273]
  PIN HI[274]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 19.000 215.650 23.000 ;
    END
  END HI[274]
  PIN HI[275]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 19.000 210.130 23.000 ;
    END
  END HI[275]
  PIN HI[276]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END HI[276]
  PIN HI[277]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END HI[277]
  PIN HI[278]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END HI[278]
  PIN HI[279]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END HI[279]
  PIN HI[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 19.000 142.050 23.000 ;
    END
  END HI[27]
  PIN HI[280]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END HI[280]
  PIN HI[281]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 19.000 6.810 23.000 ;
    END
  END HI[281]
  PIN HI[282]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 19.000 135.610 23.000 ;
    END
  END HI[282]
  PIN HI[283]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END HI[283]
  PIN HI[284]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END HI[284]
  PIN HI[285]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 10.920 300.000 11.520 ;
    END
  END HI[285]
  PIN HI[286]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 19.000 80.410 23.000 ;
    END
  END HI[286]
  PIN HI[287]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 19.000 126.410 23.000 ;
    END
  END HI[287]
  PIN HI[288]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 19.000 203.690 23.000 ;
    END
  END HI[288]
  PIN HI[289]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 19.000 110.770 23.000 ;
    END
  END HI[289]
  PIN HI[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END HI[28]
  PIN HI[290]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 19.000 199.090 23.000 ;
    END
  END HI[290]
  PIN HI[291]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 19.000 35.330 23.000 ;
    END
  END HI[291]
  PIN HI[292]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 19.000 12.330 23.000 ;
    END
  END HI[292]
  PIN HI[293]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END HI[293]
  PIN HI[294]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END HI[294]
  PIN HI[295]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END HI[295]
  PIN HI[296]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END HI[296]
  PIN HI[297]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END HI[297]
  PIN HI[298]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 19.000 268.090 23.000 ;
    END
  END HI[298]
  PIN HI[299]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END HI[299]
  PIN HI[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END HI[29]
  PIN HI[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 19.000 213.810 23.000 ;
    END
  END HI[2]
  PIN HI[300]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 19.000 73.050 23.000 ;
    END
  END HI[300]
  PIN HI[301]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END HI[301]
  PIN HI[302]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END HI[302]
  PIN HI[303]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END HI[303]
  PIN HI[304]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 19.000 54.650 23.000 ;
    END
  END HI[304]
  PIN HI[305]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END HI[305]
  PIN HI[306]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 19.000 24.290 23.000 ;
    END
  END HI[306]
  PIN HI[307]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END HI[307]
  PIN HI[308]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 19.000 53.730 23.000 ;
    END
  END HI[308]
  PIN HI[309]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 19.000 164.130 23.000 ;
    END
  END HI[309]
  PIN HI[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END HI[30]
  PIN HI[310]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END HI[310]
  PIN HI[311]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END HI[311]
  PIN HI[312]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 19.000 11.410 23.000 ;
    END
  END HI[312]
  PIN HI[313]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END HI[313]
  PIN HI[314]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END HI[314]
  PIN HI[315]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END HI[315]
  PIN HI[316]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 19.000 264.410 23.000 ;
    END
  END HI[316]
  PIN HI[317]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END HI[317]
  PIN HI[318]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END HI[318]
  PIN HI[319]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END HI[319]
  PIN HI[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END HI[31]
  PIN HI[320]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END HI[320]
  PIN HI[321]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END HI[321]
  PIN HI[322]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 19.000 288.330 23.000 ;
    END
  END HI[322]
  PIN HI[323]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END HI[323]
  PIN HI[324]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END HI[324]
  PIN HI[325]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 19.000 119.050 23.000 ;
    END
  END HI[325]
  PIN HI[326]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END HI[326]
  PIN HI[327]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END HI[327]
  PIN HI[328]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 19.000 179.770 23.000 ;
    END
  END HI[328]
  PIN HI[329]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END HI[329]
  PIN HI[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 19.000 257.970 23.000 ;
    END
  END HI[32]
  PIN HI[330]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END HI[330]
  PIN HI[331]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END HI[331]
  PIN HI[332]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 19.000 168.730 23.000 ;
    END
  END HI[332]
  PIN HI[333]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 19.000 204.610 23.000 ;
    END
  END HI[333]
  PIN HI[334]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END HI[334]
  PIN HI[335]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END HI[335]
  PIN HI[336]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 19.000 290.170 23.000 ;
    END
  END HI[336]
  PIN HI[337]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 19.000 225.770 23.000 ;
    END
  END HI[337]
  PIN HI[338]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 19.000 182.530 23.000 ;
    END
  END HI[338]
  PIN HI[339]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 19.000 56.490 23.000 ;
    END
  END HI[339]
  PIN HI[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END HI[33]
  PIN HI[340]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 19.000 162.290 23.000 ;
    END
  END HI[340]
  PIN HI[341]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END HI[341]
  PIN HI[342]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 19.000 125.490 23.000 ;
    END
  END HI[342]
  PIN HI[343]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END HI[343]
  PIN HI[344]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END HI[344]
  PIN HI[345]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END HI[345]
  PIN HI[346]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END HI[346]
  PIN HI[347]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 19.000 99.730 23.000 ;
    END
  END HI[347]
  PIN HI[348]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 19.000 119.970 23.000 ;
    END
  END HI[348]
  PIN HI[349]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END HI[349]
  PIN HI[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END HI[34]
  PIN HI[350]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 19.000 29.810 23.000 ;
    END
  END HI[350]
  PIN HI[351]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END HI[351]
  PIN HI[352]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 19.000 240.490 23.000 ;
    END
  END HI[352]
  PIN HI[353]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 19.000 83.170 23.000 ;
    END
  END HI[353]
  PIN HI[354]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 19.000 224.850 23.000 ;
    END
  END HI[354]
  PIN HI[355]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 19.000 32.570 23.000 ;
    END
  END HI[355]
  PIN HI[356]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 19.000 252.450 23.000 ;
    END
  END HI[356]
  PIN HI[357]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END HI[357]
  PIN HI[358]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 19.000 177.010 23.000 ;
    END
  END HI[358]
  PIN HI[359]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 19.000 218.410 23.000 ;
    END
  END HI[359]
  PIN HI[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 19.000 270.850 23.000 ;
    END
  END HI[35]
  PIN HI[360]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END HI[360]
  PIN HI[361]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 8.200 300.000 8.800 ;
    END
  END HI[361]
  PIN HI[362]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END HI[362]
  PIN HI[363]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 5.480 300.000 6.080 ;
    END
  END HI[363]
  PIN HI[364]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 19.000 146.650 23.000 ;
    END
  END HI[364]
  PIN HI[365]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END HI[365]
  PIN HI[366]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 19.000 140.210 23.000 ;
    END
  END HI[366]
  PIN HI[367]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END HI[367]
  PIN HI[368]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END HI[368]
  PIN HI[369]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END HI[369]
  PIN HI[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END HI[36]
  PIN HI[370]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 19.000 249.690 23.000 ;
    END
  END HI[370]
  PIN HI[371]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END HI[371]
  PIN HI[372]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 19.000 107.090 23.000 ;
    END
  END HI[372]
  PIN HI[373]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END HI[373]
  PIN HI[374]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 19.000 147.570 23.000 ;
    END
  END HI[374]
  PIN HI[375]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 19.000 132.850 23.000 ;
    END
  END HI[375]
  PIN HI[376]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 19.000 269.930 23.000 ;
    END
  END HI[376]
  PIN HI[377]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 19.000 48.210 23.000 ;
    END
  END HI[377]
  PIN HI[378]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END HI[378]
  PIN HI[379]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END HI[379]
  PIN HI[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 19.000 84.090 23.000 ;
    END
  END HI[37]
  PIN HI[380]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 19.000 192.650 23.000 ;
    END
  END HI[380]
  PIN HI[381]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 19.000 3.130 23.000 ;
    END
  END HI[381]
  PIN HI[382]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END HI[382]
  PIN HI[383]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 19.000 33.490 23.000 ;
    END
  END HI[383]
  PIN HI[384]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END HI[384]
  PIN HI[385]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 19.000 150.330 23.000 ;
    END
  END HI[385]
  PIN HI[386]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END HI[386]
  PIN HI[387]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 19.000 228.530 23.000 ;
    END
  END HI[387]
  PIN HI[388]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END HI[388]
  PIN HI[389]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 19.000 159.530 23.000 ;
    END
  END HI[389]
  PIN HI[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 19.000 116.290 23.000 ;
    END
  END HI[38]
  PIN HI[390]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END HI[390]
  PIN HI[391]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END HI[391]
  PIN HI[392]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END HI[392]
  PIN HI[393]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 19.000 237.730 23.000 ;
    END
  END HI[393]
  PIN HI[394]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END HI[394]
  PIN HI[395]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 19.000 105.250 23.000 ;
    END
  END HI[395]
  PIN HI[396]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 19.000 285.570 23.000 ;
    END
  END HI[396]
  PIN HI[397]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END HI[397]
  PIN HI[398]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 19.000 143.890 23.000 ;
    END
  END HI[398]
  PIN HI[399]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 19.000 114.450 23.000 ;
    END
  END HI[399]
  PIN HI[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END HI[39]
  PIN HI[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END HI[3]
  PIN HI[400]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END HI[400]
  PIN HI[401]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END HI[401]
  PIN HI[402]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 19.000 78.570 23.000 ;
    END
  END HI[402]
  PIN HI[403]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 19.000 38.090 23.000 ;
    END
  END HI[403]
  PIN HI[404]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 19.000 282.810 23.000 ;
    END
  END HI[404]
  PIN HI[405]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END HI[405]
  PIN HI[406]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END HI[406]
  PIN HI[407]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END HI[407]
  PIN HI[408]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 19.000 44.530 23.000 ;
    END
  END HI[408]
  PIN HI[409]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 19.000 188.050 23.000 ;
    END
  END HI[409]
  PIN HI[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END HI[40]
  PIN HI[410]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END HI[410]
  PIN HI[411]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END HI[411]
  PIN HI[412]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END HI[412]
  PIN HI[413]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END HI[413]
  PIN HI[414]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END HI[414]
  PIN HI[415]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END HI[415]
  PIN HI[416]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 19.000 152.170 23.000 ;
    END
  END HI[416]
  PIN HI[417]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END HI[417]
  PIN HI[418]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 19.000 279.130 23.000 ;
    END
  END HI[418]
  PIN HI[419]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END HI[419]
  PIN HI[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 19.000 171.490 23.000 ;
    END
  END HI[41]
  PIN HI[420]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END HI[420]
  PIN HI[421]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 19.000 75.810 23.000 ;
    END
  END HI[421]
  PIN HI[422]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 19.000 60.170 23.000 ;
    END
  END HI[422]
  PIN HI[423]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END HI[423]
  PIN HI[424]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END HI[424]
  PIN HI[425]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 19.000 291.090 23.000 ;
    END
  END HI[425]
  PIN HI[426]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 19.000 50.050 23.000 ;
    END
  END HI[426]
  PIN HI[427]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 19.000 293.850 23.000 ;
    END
  END HI[427]
  PIN HI[428]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END HI[428]
  PIN HI[429]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END HI[429]
  PIN HI[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END HI[42]
  PIN HI[430]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 19.000 180.690 23.000 ;
    END
  END HI[430]
  PIN HI[431]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 19.000 173.330 23.000 ;
    END
  END HI[431]
  PIN HI[432]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 19.000 86.850 23.000 ;
    END
  END HI[432]
  PIN HI[433]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 19.000 90.530 23.000 ;
    END
  END HI[433]
  PIN HI[434]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 19.000 242.330 23.000 ;
    END
  END HI[434]
  PIN HI[435]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 19.000 81.330 23.000 ;
    END
  END HI[435]
  PIN HI[436]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END HI[436]
  PIN HI[437]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END HI[437]
  PIN HI[438]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 19.000 275.450 23.000 ;
    END
  END HI[438]
  PIN HI[439]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 13.640 300.000 14.240 ;
    END
  END HI[439]
  PIN HI[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END HI[43]
  PIN HI[440]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END HI[440]
  PIN HI[441]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 19.000 234.050 23.000 ;
    END
  END HI[441]
  PIN HI[442]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 19.000 69.370 23.000 ;
    END
  END HI[442]
  PIN HI[443]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 19.000 260.730 23.000 ;
    END
  END HI[443]
  PIN HI[444]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 19.000 71.210 23.000 ;
    END
  END HI[444]
  PIN HI[445]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 19.000 129.170 23.000 ;
    END
  END HI[445]
  PIN HI[446]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END HI[446]
  PIN HI[447]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END HI[447]
  PIN HI[448]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END HI[448]
  PIN HI[449]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END HI[449]
  PIN HI[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 19.000 41.770 23.000 ;
    END
  END HI[44]
  PIN HI[450]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 19.000 92.370 23.000 ;
    END
  END HI[450]
  PIN HI[451]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END HI[451]
  PIN HI[452]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END HI[452]
  PIN HI[453]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 19.000 27.970 23.000 ;
    END
  END HI[453]
  PIN HI[454]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 19.000 122.730 23.000 ;
    END
  END HI[454]
  PIN HI[455]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END HI[455]
  PIN HI[456]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END HI[456]
  PIN HI[457]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 19.000 89.610 23.000 ;
    END
  END HI[457]
  PIN HI[458]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END HI[458]
  PIN HI[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 19.000 201.850 23.000 ;
    END
  END HI[45]
  PIN HI[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END HI[46]
  PIN HI[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END HI[47]
  PIN HI[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END HI[48]
  PIN HI[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 19.000 154.010 23.000 ;
    END
  END HI[49]
  PIN HI[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END HI[4]
  PIN HI[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END HI[50]
  PIN HI[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END HI[51]
  PIN HI[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 19.000 245.090 23.000 ;
    END
  END HI[52]
  PIN HI[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 19.000 101.570 23.000 ;
    END
  END HI[53]
  PIN HI[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 19.000 287.410 23.000 ;
    END
  END HI[54]
  PIN HI[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END HI[55]
  PIN HI[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END HI[56]
  PIN HI[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 19.000 280.050 23.000 ;
    END
  END HI[57]
  PIN HI[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 19.000 96.970 23.000 ;
    END
  END HI[58]
  PIN HI[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END HI[59]
  PIN HI[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 19.000 176.090 23.000 ;
    END
  END HI[5]
  PIN HI[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 19.000 251.530 23.000 ;
    END
  END HI[60]
  PIN HI[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END HI[61]
  PIN HI[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END HI[62]
  PIN HI[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END HI[63]
  PIN HI[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END HI[64]
  PIN HI[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END HI[65]
  PIN HI[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END HI[66]
  PIN HI[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END HI[67]
  PIN HI[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END HI[68]
  PIN HI[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END HI[69]
  PIN HI[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END HI[6]
  PIN HI[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 19.000 17.850 23.000 ;
    END
  END HI[70]
  PIN HI[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END HI[71]
  PIN HI[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 19.000 20.610 23.000 ;
    END
  END HI[72]
  PIN HI[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 19.000 68.450 23.000 ;
    END
  END HI[73]
  PIN HI[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END HI[74]
  PIN HI[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 19.000 248.770 23.000 ;
    END
  END HI[75]
  PIN HI[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 19.000 223.010 23.000 ;
    END
  END HI[76]
  PIN HI[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 19.000 167.810 23.000 ;
    END
  END HI[77]
  PIN HI[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 19.000 246.010 23.000 ;
    END
  END HI[78]
  PIN HI[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 19.000 233.130 23.000 ;
    END
  END HI[79]
  PIN HI[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END HI[7]
  PIN HI[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 19.000 161.370 23.000 ;
    END
  END HI[80]
  PIN HI[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 19.000 257.050 23.000 ;
    END
  END HI[81]
  PIN HI[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END HI[82]
  PIN HI[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 19.000 87.770 23.000 ;
    END
  END HI[83]
  PIN HI[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 19.000 104.330 23.000 ;
    END
  END HI[84]
  PIN HI[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 19.000 50.970 23.000 ;
    END
  END HI[85]
  PIN HI[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 19.000 155.850 23.000 ;
    END
  END HI[86]
  PIN HI[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END HI[87]
  PIN HI[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 19.000 266.250 23.000 ;
    END
  END HI[88]
  PIN HI[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 19.000 9.570 23.000 ;
    END
  END HI[89]
  PIN HI[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 19.000 189.890 23.000 ;
    END
  END HI[8]
  PIN HI[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 19.000 5.890 23.000 ;
    END
  END HI[90]
  PIN HI[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 19.000 134.690 23.000 ;
    END
  END HI[91]
  PIN HI[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 19.000 16.010 23.000 ;
    END
  END HI[92]
  PIN HI[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END HI[93]
  PIN HI[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 19.000 230.370 23.000 ;
    END
  END HI[94]
  PIN HI[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 19.000 14.170 23.000 ;
    END
  END HI[95]
  PIN HI[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END HI[96]
  PIN HI[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 19.000 77.650 23.000 ;
    END
  END HI[97]
  PIN HI[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END HI[98]
  PIN HI[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 4.120 300.000 4.720 ;
    END
  END HI[99]
  PIN HI[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END HI[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 256.750 5.200 257.050 16.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 176.750 5.200 177.050 16.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 96.750 5.200 97.050 16.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 16.750 5.200 17.050 16.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 6.900 6.050 293.020 6.350 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 216.750 5.200 217.050 16.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 136.750 5.200 137.050 16.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 56.750 5.200 57.050 16.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 6.900 11.450 293.020 11.750 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 6.900 5.355 293.020 16.405 ;
      LAYER met1 ;
        RECT 2.830 4.460 296.630 17.640 ;
      LAYER met2 ;
        RECT 3.410 18.720 3.490 19.000 ;
        RECT 4.330 18.720 5.330 19.000 ;
        RECT 6.170 18.720 6.250 19.000 ;
        RECT 7.090 18.720 8.090 19.000 ;
        RECT 8.930 18.720 9.010 19.000 ;
        RECT 9.850 18.720 10.850 19.000 ;
        RECT 11.690 18.720 11.770 19.000 ;
        RECT 12.610 18.720 13.610 19.000 ;
        RECT 14.450 18.720 14.530 19.000 ;
        RECT 15.370 18.720 15.450 19.000 ;
        RECT 16.290 18.720 17.290 19.000 ;
        RECT 18.130 18.720 18.210 19.000 ;
        RECT 19.050 18.720 20.050 19.000 ;
        RECT 20.890 18.720 20.970 19.000 ;
        RECT 21.810 18.720 22.810 19.000 ;
        RECT 23.650 18.720 23.730 19.000 ;
        RECT 24.570 18.720 25.570 19.000 ;
        RECT 26.410 18.720 26.490 19.000 ;
        RECT 27.330 18.720 27.410 19.000 ;
        RECT 28.250 18.720 29.250 19.000 ;
        RECT 30.090 18.720 30.170 19.000 ;
        RECT 31.010 18.720 32.010 19.000 ;
        RECT 32.850 18.720 32.930 19.000 ;
        RECT 33.770 18.720 34.770 19.000 ;
        RECT 35.610 18.720 35.690 19.000 ;
        RECT 36.530 18.720 37.530 19.000 ;
        RECT 38.370 18.720 38.450 19.000 ;
        RECT 39.290 18.720 39.370 19.000 ;
        RECT 40.210 18.720 41.210 19.000 ;
        RECT 42.050 18.720 42.130 19.000 ;
        RECT 42.970 18.720 43.970 19.000 ;
        RECT 44.810 18.720 44.890 19.000 ;
        RECT 45.730 18.720 46.730 19.000 ;
        RECT 47.570 18.720 47.650 19.000 ;
        RECT 48.490 18.720 49.490 19.000 ;
        RECT 50.330 18.720 50.410 19.000 ;
        RECT 51.250 18.720 51.330 19.000 ;
        RECT 52.170 18.720 53.170 19.000 ;
        RECT 54.010 18.720 54.090 19.000 ;
        RECT 54.930 18.720 55.930 19.000 ;
        RECT 56.770 18.720 56.850 19.000 ;
        RECT 57.690 18.720 58.690 19.000 ;
        RECT 59.530 18.720 59.610 19.000 ;
        RECT 60.450 18.720 60.530 19.000 ;
        RECT 61.370 18.720 62.370 19.000 ;
        RECT 63.210 18.720 63.290 19.000 ;
        RECT 64.130 18.720 65.130 19.000 ;
        RECT 65.970 18.720 66.050 19.000 ;
        RECT 66.890 18.720 67.890 19.000 ;
        RECT 68.730 18.720 68.810 19.000 ;
        RECT 69.650 18.720 70.650 19.000 ;
        RECT 71.490 18.720 71.570 19.000 ;
        RECT 72.410 18.720 72.490 19.000 ;
        RECT 73.330 18.720 74.330 19.000 ;
        RECT 75.170 18.720 75.250 19.000 ;
        RECT 76.090 18.720 77.090 19.000 ;
        RECT 77.930 18.720 78.010 19.000 ;
        RECT 78.850 18.720 79.850 19.000 ;
        RECT 80.690 18.720 80.770 19.000 ;
        RECT 81.610 18.720 82.610 19.000 ;
        RECT 83.450 18.720 83.530 19.000 ;
        RECT 84.370 18.720 84.450 19.000 ;
        RECT 85.290 18.720 86.290 19.000 ;
        RECT 87.130 18.720 87.210 19.000 ;
        RECT 88.050 18.720 89.050 19.000 ;
        RECT 89.890 18.720 89.970 19.000 ;
        RECT 90.810 18.720 91.810 19.000 ;
        RECT 92.650 18.720 92.730 19.000 ;
        RECT 93.570 18.720 94.570 19.000 ;
        RECT 95.410 18.720 95.490 19.000 ;
        RECT 96.330 18.720 96.410 19.000 ;
        RECT 97.250 18.720 98.250 19.000 ;
        RECT 99.090 18.720 99.170 19.000 ;
        RECT 100.010 18.720 101.010 19.000 ;
        RECT 101.850 18.720 101.930 19.000 ;
        RECT 102.770 18.720 103.770 19.000 ;
        RECT 104.610 18.720 104.690 19.000 ;
        RECT 105.530 18.720 106.530 19.000 ;
        RECT 107.370 18.720 107.450 19.000 ;
        RECT 108.290 18.720 108.370 19.000 ;
        RECT 109.210 18.720 110.210 19.000 ;
        RECT 111.050 18.720 111.130 19.000 ;
        RECT 111.970 18.720 112.970 19.000 ;
        RECT 113.810 18.720 113.890 19.000 ;
        RECT 114.730 18.720 115.730 19.000 ;
        RECT 116.570 18.720 116.650 19.000 ;
        RECT 117.490 18.720 118.490 19.000 ;
        RECT 119.330 18.720 119.410 19.000 ;
        RECT 120.250 18.720 120.330 19.000 ;
        RECT 121.170 18.720 122.170 19.000 ;
        RECT 123.010 18.720 123.090 19.000 ;
        RECT 123.930 18.720 124.930 19.000 ;
        RECT 125.770 18.720 125.850 19.000 ;
        RECT 126.690 18.720 127.690 19.000 ;
        RECT 128.530 18.720 128.610 19.000 ;
        RECT 129.450 18.720 129.530 19.000 ;
        RECT 130.370 18.720 131.370 19.000 ;
        RECT 132.210 18.720 132.290 19.000 ;
        RECT 133.130 18.720 134.130 19.000 ;
        RECT 134.970 18.720 135.050 19.000 ;
        RECT 135.890 18.720 136.890 19.000 ;
        RECT 137.730 18.720 137.810 19.000 ;
        RECT 138.650 18.720 139.650 19.000 ;
        RECT 140.490 18.720 140.570 19.000 ;
        RECT 141.410 18.720 141.490 19.000 ;
        RECT 142.330 18.720 143.330 19.000 ;
        RECT 144.170 18.720 144.250 19.000 ;
        RECT 145.090 18.720 146.090 19.000 ;
        RECT 146.930 18.720 147.010 19.000 ;
        RECT 147.850 18.720 148.850 19.000 ;
        RECT 149.690 18.720 149.770 19.000 ;
        RECT 150.610 18.720 151.610 19.000 ;
        RECT 152.450 18.720 152.530 19.000 ;
        RECT 153.370 18.720 153.450 19.000 ;
        RECT 154.290 18.720 155.290 19.000 ;
        RECT 156.130 18.720 156.210 19.000 ;
        RECT 157.050 18.720 158.050 19.000 ;
        RECT 158.890 18.720 158.970 19.000 ;
        RECT 159.810 18.720 160.810 19.000 ;
        RECT 161.650 18.720 161.730 19.000 ;
        RECT 162.570 18.720 163.570 19.000 ;
        RECT 164.410 18.720 164.490 19.000 ;
        RECT 165.330 18.720 165.410 19.000 ;
        RECT 166.250 18.720 167.250 19.000 ;
        RECT 168.090 18.720 168.170 19.000 ;
        RECT 169.010 18.720 170.010 19.000 ;
        RECT 170.850 18.720 170.930 19.000 ;
        RECT 171.770 18.720 172.770 19.000 ;
        RECT 173.610 18.720 173.690 19.000 ;
        RECT 174.530 18.720 175.530 19.000 ;
        RECT 176.370 18.720 176.450 19.000 ;
        RECT 177.290 18.720 177.370 19.000 ;
        RECT 178.210 18.720 179.210 19.000 ;
        RECT 180.050 18.720 180.130 19.000 ;
        RECT 180.970 18.720 181.970 19.000 ;
        RECT 182.810 18.720 182.890 19.000 ;
        RECT 183.730 18.720 184.730 19.000 ;
        RECT 185.570 18.720 185.650 19.000 ;
        RECT 186.490 18.720 187.490 19.000 ;
        RECT 188.330 18.720 188.410 19.000 ;
        RECT 189.250 18.720 189.330 19.000 ;
        RECT 190.170 18.720 191.170 19.000 ;
        RECT 192.010 18.720 192.090 19.000 ;
        RECT 192.930 18.720 193.930 19.000 ;
        RECT 194.770 18.720 194.850 19.000 ;
        RECT 195.690 18.720 196.690 19.000 ;
        RECT 197.530 18.720 197.610 19.000 ;
        RECT 198.450 18.720 198.530 19.000 ;
        RECT 199.370 18.720 200.370 19.000 ;
        RECT 201.210 18.720 201.290 19.000 ;
        RECT 202.130 18.720 203.130 19.000 ;
        RECT 203.970 18.720 204.050 19.000 ;
        RECT 204.890 18.720 205.890 19.000 ;
        RECT 206.730 18.720 206.810 19.000 ;
        RECT 207.650 18.720 208.650 19.000 ;
        RECT 209.490 18.720 209.570 19.000 ;
        RECT 210.410 18.720 210.490 19.000 ;
        RECT 211.330 18.720 212.330 19.000 ;
        RECT 213.170 18.720 213.250 19.000 ;
        RECT 214.090 18.720 215.090 19.000 ;
        RECT 215.930 18.720 216.010 19.000 ;
        RECT 216.850 18.720 217.850 19.000 ;
        RECT 218.690 18.720 218.770 19.000 ;
        RECT 219.610 18.720 220.610 19.000 ;
        RECT 221.450 18.720 221.530 19.000 ;
        RECT 222.370 18.720 222.450 19.000 ;
        RECT 223.290 18.720 224.290 19.000 ;
        RECT 225.130 18.720 225.210 19.000 ;
        RECT 226.050 18.720 227.050 19.000 ;
        RECT 227.890 18.720 227.970 19.000 ;
        RECT 228.810 18.720 229.810 19.000 ;
        RECT 230.650 18.720 230.730 19.000 ;
        RECT 231.570 18.720 232.570 19.000 ;
        RECT 233.410 18.720 233.490 19.000 ;
        RECT 234.330 18.720 234.410 19.000 ;
        RECT 235.250 18.720 236.250 19.000 ;
        RECT 237.090 18.720 237.170 19.000 ;
        RECT 238.010 18.720 239.010 19.000 ;
        RECT 239.850 18.720 239.930 19.000 ;
        RECT 240.770 18.720 241.770 19.000 ;
        RECT 242.610 18.720 242.690 19.000 ;
        RECT 243.530 18.720 244.530 19.000 ;
        RECT 245.370 18.720 245.450 19.000 ;
        RECT 246.290 18.720 246.370 19.000 ;
        RECT 247.210 18.720 248.210 19.000 ;
        RECT 249.050 18.720 249.130 19.000 ;
        RECT 249.970 18.720 250.970 19.000 ;
        RECT 251.810 18.720 251.890 19.000 ;
        RECT 252.730 18.720 253.730 19.000 ;
        RECT 254.570 18.720 254.650 19.000 ;
        RECT 255.490 18.720 256.490 19.000 ;
        RECT 257.330 18.720 257.410 19.000 ;
        RECT 258.250 18.720 258.330 19.000 ;
        RECT 259.170 18.720 260.170 19.000 ;
        RECT 261.010 18.720 261.090 19.000 ;
        RECT 261.930 18.720 262.930 19.000 ;
        RECT 263.770 18.720 263.850 19.000 ;
        RECT 264.690 18.720 265.690 19.000 ;
        RECT 266.530 18.720 266.610 19.000 ;
        RECT 267.450 18.720 267.530 19.000 ;
        RECT 268.370 18.720 269.370 19.000 ;
        RECT 270.210 18.720 270.290 19.000 ;
        RECT 271.130 18.720 272.130 19.000 ;
        RECT 272.970 18.720 273.050 19.000 ;
        RECT 273.890 18.720 274.890 19.000 ;
        RECT 275.730 18.720 275.810 19.000 ;
        RECT 276.650 18.720 277.650 19.000 ;
        RECT 278.490 18.720 278.570 19.000 ;
        RECT 279.410 18.720 279.490 19.000 ;
        RECT 280.330 18.720 281.330 19.000 ;
        RECT 282.170 18.720 282.250 19.000 ;
        RECT 283.090 18.720 284.090 19.000 ;
        RECT 284.930 18.720 285.010 19.000 ;
        RECT 285.850 18.720 286.850 19.000 ;
        RECT 287.690 18.720 287.770 19.000 ;
        RECT 288.610 18.720 289.610 19.000 ;
        RECT 290.450 18.720 290.530 19.000 ;
        RECT 291.370 18.720 291.450 19.000 ;
        RECT 292.290 18.720 293.290 19.000 ;
        RECT 294.130 18.720 294.210 19.000 ;
        RECT 295.050 18.720 296.050 19.000 ;
        RECT 2.860 16.840 296.600 18.720 ;
        RECT 2.860 4.920 16.470 16.840 ;
        RECT 17.330 4.920 56.470 16.840 ;
        RECT 57.330 4.920 96.470 16.840 ;
        RECT 97.330 4.920 136.470 16.840 ;
        RECT 137.330 4.920 176.470 16.840 ;
        RECT 177.330 4.920 216.470 16.840 ;
        RECT 217.330 4.920 256.470 16.840 ;
        RECT 257.330 4.920 296.600 16.840 ;
        RECT 2.860 4.280 296.600 4.920 ;
        RECT 3.410 0.155 3.490 4.280 ;
        RECT 4.330 0.155 4.410 4.280 ;
        RECT 5.250 0.155 6.250 4.280 ;
        RECT 7.090 0.155 7.170 4.280 ;
        RECT 8.010 0.155 9.010 4.280 ;
        RECT 9.850 0.155 9.930 4.280 ;
        RECT 10.770 0.155 11.770 4.280 ;
        RECT 12.610 0.155 12.690 4.280 ;
        RECT 13.530 0.155 13.610 4.280 ;
        RECT 14.450 0.155 15.450 4.280 ;
        RECT 16.290 0.155 16.370 4.280 ;
        RECT 17.210 0.155 18.210 4.280 ;
        RECT 19.050 0.155 19.130 4.280 ;
        RECT 19.970 0.155 20.970 4.280 ;
        RECT 21.810 0.155 21.890 4.280 ;
        RECT 22.730 0.155 23.730 4.280 ;
        RECT 24.570 0.155 24.650 4.280 ;
        RECT 25.490 0.155 25.570 4.280 ;
        RECT 26.410 0.155 27.410 4.280 ;
        RECT 28.250 0.155 28.330 4.280 ;
        RECT 29.170 0.155 30.170 4.280 ;
        RECT 31.010 0.155 31.090 4.280 ;
        RECT 31.930 0.155 32.930 4.280 ;
        RECT 33.770 0.155 33.850 4.280 ;
        RECT 34.690 0.155 35.690 4.280 ;
        RECT 36.530 0.155 36.610 4.280 ;
        RECT 37.450 0.155 37.530 4.280 ;
        RECT 38.370 0.155 39.370 4.280 ;
        RECT 40.210 0.155 40.290 4.280 ;
        RECT 41.130 0.155 42.130 4.280 ;
        RECT 42.970 0.155 43.050 4.280 ;
        RECT 43.890 0.155 44.890 4.280 ;
        RECT 45.730 0.155 45.810 4.280 ;
        RECT 46.650 0.155 47.650 4.280 ;
        RECT 48.490 0.155 48.570 4.280 ;
        RECT 49.410 0.155 49.490 4.280 ;
        RECT 50.330 0.155 51.330 4.280 ;
        RECT 52.170 0.155 52.250 4.280 ;
        RECT 53.090 0.155 54.090 4.280 ;
        RECT 54.930 0.155 55.010 4.280 ;
        RECT 55.850 0.155 56.850 4.280 ;
        RECT 57.690 0.155 57.770 4.280 ;
        RECT 58.610 0.155 59.610 4.280 ;
        RECT 60.450 0.155 60.530 4.280 ;
        RECT 61.370 0.155 61.450 4.280 ;
        RECT 62.290 0.155 63.290 4.280 ;
        RECT 64.130 0.155 64.210 4.280 ;
        RECT 65.050 0.155 66.050 4.280 ;
        RECT 66.890 0.155 66.970 4.280 ;
        RECT 67.810 0.155 68.810 4.280 ;
        RECT 69.650 0.155 69.730 4.280 ;
        RECT 70.570 0.155 70.650 4.280 ;
        RECT 71.490 0.155 72.490 4.280 ;
        RECT 73.330 0.155 73.410 4.280 ;
        RECT 74.250 0.155 75.250 4.280 ;
        RECT 76.090 0.155 76.170 4.280 ;
        RECT 77.010 0.155 78.010 4.280 ;
        RECT 78.850 0.155 78.930 4.280 ;
        RECT 79.770 0.155 80.770 4.280 ;
        RECT 81.610 0.155 81.690 4.280 ;
        RECT 82.530 0.155 82.610 4.280 ;
        RECT 83.450 0.155 84.450 4.280 ;
        RECT 85.290 0.155 85.370 4.280 ;
        RECT 86.210 0.155 87.210 4.280 ;
        RECT 88.050 0.155 88.130 4.280 ;
        RECT 88.970 0.155 89.970 4.280 ;
        RECT 90.810 0.155 90.890 4.280 ;
        RECT 91.730 0.155 92.730 4.280 ;
        RECT 93.570 0.155 93.650 4.280 ;
        RECT 94.490 0.155 94.570 4.280 ;
        RECT 95.410 0.155 96.410 4.280 ;
        RECT 97.250 0.155 97.330 4.280 ;
        RECT 98.170 0.155 99.170 4.280 ;
        RECT 100.010 0.155 100.090 4.280 ;
        RECT 100.930 0.155 101.930 4.280 ;
        RECT 102.770 0.155 102.850 4.280 ;
        RECT 103.690 0.155 104.690 4.280 ;
        RECT 105.530 0.155 105.610 4.280 ;
        RECT 106.450 0.155 106.530 4.280 ;
        RECT 107.370 0.155 108.370 4.280 ;
        RECT 109.210 0.155 109.290 4.280 ;
        RECT 110.130 0.155 111.130 4.280 ;
        RECT 111.970 0.155 112.050 4.280 ;
        RECT 112.890 0.155 113.890 4.280 ;
        RECT 114.730 0.155 114.810 4.280 ;
        RECT 115.650 0.155 116.650 4.280 ;
        RECT 117.490 0.155 117.570 4.280 ;
        RECT 118.410 0.155 118.490 4.280 ;
        RECT 119.330 0.155 120.330 4.280 ;
        RECT 121.170 0.155 121.250 4.280 ;
        RECT 122.090 0.155 123.090 4.280 ;
        RECT 123.930 0.155 124.010 4.280 ;
        RECT 124.850 0.155 125.850 4.280 ;
        RECT 126.690 0.155 126.770 4.280 ;
        RECT 127.610 0.155 128.610 4.280 ;
        RECT 129.450 0.155 129.530 4.280 ;
        RECT 130.370 0.155 130.450 4.280 ;
        RECT 131.290 0.155 132.290 4.280 ;
        RECT 133.130 0.155 133.210 4.280 ;
        RECT 134.050 0.155 135.050 4.280 ;
        RECT 135.890 0.155 135.970 4.280 ;
        RECT 136.810 0.155 137.810 4.280 ;
        RECT 138.650 0.155 138.730 4.280 ;
        RECT 139.570 0.155 139.650 4.280 ;
        RECT 140.490 0.155 141.490 4.280 ;
        RECT 142.330 0.155 142.410 4.280 ;
        RECT 143.250 0.155 144.250 4.280 ;
        RECT 145.090 0.155 145.170 4.280 ;
        RECT 146.010 0.155 147.010 4.280 ;
        RECT 147.850 0.155 147.930 4.280 ;
        RECT 148.770 0.155 149.770 4.280 ;
        RECT 150.610 0.155 150.690 4.280 ;
        RECT 151.530 0.155 151.610 4.280 ;
        RECT 152.450 0.155 153.450 4.280 ;
        RECT 154.290 0.155 154.370 4.280 ;
        RECT 155.210 0.155 156.210 4.280 ;
        RECT 157.050 0.155 157.130 4.280 ;
        RECT 157.970 0.155 158.970 4.280 ;
        RECT 159.810 0.155 159.890 4.280 ;
        RECT 160.730 0.155 161.730 4.280 ;
        RECT 162.570 0.155 162.650 4.280 ;
        RECT 163.490 0.155 163.570 4.280 ;
        RECT 164.410 0.155 165.410 4.280 ;
        RECT 166.250 0.155 166.330 4.280 ;
        RECT 167.170 0.155 168.170 4.280 ;
        RECT 169.010 0.155 169.090 4.280 ;
        RECT 169.930 0.155 170.930 4.280 ;
        RECT 171.770 0.155 171.850 4.280 ;
        RECT 172.690 0.155 173.690 4.280 ;
        RECT 174.530 0.155 174.610 4.280 ;
        RECT 175.450 0.155 175.530 4.280 ;
        RECT 176.370 0.155 177.370 4.280 ;
        RECT 178.210 0.155 178.290 4.280 ;
        RECT 179.130 0.155 180.130 4.280 ;
        RECT 180.970 0.155 181.050 4.280 ;
        RECT 181.890 0.155 182.890 4.280 ;
        RECT 183.730 0.155 183.810 4.280 ;
        RECT 184.650 0.155 185.650 4.280 ;
        RECT 186.490 0.155 186.570 4.280 ;
        RECT 187.410 0.155 187.490 4.280 ;
        RECT 188.330 0.155 189.330 4.280 ;
        RECT 190.170 0.155 190.250 4.280 ;
        RECT 191.090 0.155 192.090 4.280 ;
        RECT 192.930 0.155 193.010 4.280 ;
        RECT 193.850 0.155 194.850 4.280 ;
        RECT 195.690 0.155 195.770 4.280 ;
        RECT 196.610 0.155 197.610 4.280 ;
        RECT 198.450 0.155 198.530 4.280 ;
        RECT 199.370 0.155 199.450 4.280 ;
        RECT 200.290 0.155 201.290 4.280 ;
        RECT 202.130 0.155 202.210 4.280 ;
        RECT 203.050 0.155 204.050 4.280 ;
        RECT 204.890 0.155 204.970 4.280 ;
        RECT 205.810 0.155 206.810 4.280 ;
        RECT 207.650 0.155 207.730 4.280 ;
        RECT 208.570 0.155 208.650 4.280 ;
        RECT 209.490 0.155 210.490 4.280 ;
        RECT 211.330 0.155 211.410 4.280 ;
        RECT 212.250 0.155 213.250 4.280 ;
        RECT 214.090 0.155 214.170 4.280 ;
        RECT 215.010 0.155 216.010 4.280 ;
        RECT 216.850 0.155 216.930 4.280 ;
        RECT 217.770 0.155 218.770 4.280 ;
        RECT 219.610 0.155 219.690 4.280 ;
        RECT 220.530 0.155 220.610 4.280 ;
        RECT 221.450 0.155 222.450 4.280 ;
        RECT 223.290 0.155 223.370 4.280 ;
        RECT 224.210 0.155 225.210 4.280 ;
        RECT 226.050 0.155 226.130 4.280 ;
        RECT 226.970 0.155 227.970 4.280 ;
        RECT 228.810 0.155 228.890 4.280 ;
        RECT 229.730 0.155 230.730 4.280 ;
        RECT 231.570 0.155 231.650 4.280 ;
        RECT 232.490 0.155 232.570 4.280 ;
        RECT 233.410 0.155 234.410 4.280 ;
        RECT 235.250 0.155 235.330 4.280 ;
        RECT 236.170 0.155 237.170 4.280 ;
        RECT 238.010 0.155 238.090 4.280 ;
        RECT 238.930 0.155 239.930 4.280 ;
        RECT 240.770 0.155 240.850 4.280 ;
        RECT 241.690 0.155 242.690 4.280 ;
        RECT 243.530 0.155 243.610 4.280 ;
        RECT 244.450 0.155 244.530 4.280 ;
        RECT 245.370 0.155 246.370 4.280 ;
        RECT 247.210 0.155 247.290 4.280 ;
        RECT 248.130 0.155 249.130 4.280 ;
        RECT 249.970 0.155 250.050 4.280 ;
        RECT 250.890 0.155 251.890 4.280 ;
        RECT 252.730 0.155 252.810 4.280 ;
        RECT 253.650 0.155 254.650 4.280 ;
        RECT 255.490 0.155 255.570 4.280 ;
        RECT 256.410 0.155 256.490 4.280 ;
        RECT 257.330 0.155 258.330 4.280 ;
        RECT 259.170 0.155 259.250 4.280 ;
        RECT 260.090 0.155 261.090 4.280 ;
        RECT 261.930 0.155 262.010 4.280 ;
        RECT 262.850 0.155 263.850 4.280 ;
        RECT 264.690 0.155 264.770 4.280 ;
        RECT 265.610 0.155 266.610 4.280 ;
        RECT 267.450 0.155 267.530 4.280 ;
        RECT 268.370 0.155 268.450 4.280 ;
        RECT 269.290 0.155 270.290 4.280 ;
        RECT 271.130 0.155 271.210 4.280 ;
        RECT 272.050 0.155 273.050 4.280 ;
        RECT 273.890 0.155 273.970 4.280 ;
        RECT 274.810 0.155 275.810 4.280 ;
        RECT 276.650 0.155 276.730 4.280 ;
        RECT 277.570 0.155 277.650 4.280 ;
        RECT 278.490 0.155 279.490 4.280 ;
        RECT 280.330 0.155 280.410 4.280 ;
        RECT 281.250 0.155 282.250 4.280 ;
        RECT 283.090 0.155 283.170 4.280 ;
        RECT 284.010 0.155 285.010 4.280 ;
        RECT 285.850 0.155 285.930 4.280 ;
        RECT 286.770 0.155 287.770 4.280 ;
        RECT 288.610 0.155 288.690 4.280 ;
        RECT 289.530 0.155 289.610 4.280 ;
        RECT 290.450 0.155 291.450 4.280 ;
        RECT 292.290 0.155 292.370 4.280 ;
        RECT 293.210 0.155 294.210 4.280 ;
        RECT 295.050 0.155 295.130 4.280 ;
        RECT 295.970 0.155 296.600 4.280 ;
      LAYER met3 ;
        RECT 4.400 17.320 295.600 18.185 ;
        RECT 4.000 16.000 296.000 17.320 ;
        RECT 4.400 13.240 295.600 16.000 ;
        RECT 4.000 12.150 296.000 13.240 ;
        RECT 4.000 11.920 6.500 12.150 ;
        RECT 4.400 11.050 6.500 11.920 ;
        RECT 293.420 11.920 296.000 12.150 ;
        RECT 293.420 11.050 295.600 11.920 ;
        RECT 4.400 9.160 295.600 11.050 ;
        RECT 4.000 7.840 295.600 9.160 ;
        RECT 4.400 7.800 295.600 7.840 ;
        RECT 4.400 6.750 296.000 7.800 ;
        RECT 4.400 5.650 6.500 6.750 ;
        RECT 293.420 6.480 296.000 6.750 ;
        RECT 293.420 5.650 295.600 6.480 ;
        RECT 4.400 5.080 295.600 5.650 ;
        RECT 4.000 3.720 295.600 5.080 ;
        RECT 4.000 0.175 296.000 3.720 ;
  END
END mprj_logic_high
END LIBRARY

